library verilog;
use verilog.vl_types.all;
entity simulacao_tb is
end simulacao_tb;
